package shared_pkg; 
bit test_finished;  // signal refer to the end of the testbench
int error_count,correct_count; 
event trigger;
endpackage 